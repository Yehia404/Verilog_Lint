module adder (X, Y, S);
input    X;
input     Y;
output      S;

assign S = X * Y;
endmodule
