module adder (X, Y,S);
input X,Y;
output S;

assign S= X+Y;
endmodule



